module Random_Generator_12bits(CLK,RESET,SEED,RANDOM_RESULT);
	input CLK;
	input RESET;
	input [11:0]SEED;
	output reg [11:0]RANDOM_RESULT;

	always @(posedge CLK)begin
		if(RESET)begin
			RANDOM_RESULT<=SEED;
		end
		else begin
			RANDOM_RESULT[0]<=RANDOM_RESULT[11];
			RANDOM_RESULT[1]<=RANDOM_RESULT[0]^RANDOM_RESULT[11];
			RANDOM_RESULT[2]<=RANDOM_RESULT[1];
			RANDOM_RESULT[3]<=RANDOM_RESULT[2];
			RANDOM_RESULT[4]<=RANDOM_RESULT[3]^RANDOM_RESULT[11];
			RANDOM_RESULT[5]<=RANDOM_RESULT[4];
			RANDOM_RESULT[6]<=RANDOM_RESULT[5];
			RANDOM_RESULT[7]<=RANDOM_RESULT[6]^RANDOM_RESULT[11];
			RANDOM_RESULT[8]<=RANDOM_RESULT[7];
			RANDOM_RESULT[9]<=RANDOM_RESULT[8];
			RANDOM_RESULT[10]<=RANDOM_RESULT[9];
			RANDOM_RESULT[11]<=RANDOM_RESULT[10];
		end
	end
endmodule