module Random_Generator_16bits(CLK,RESET,SEED,RANDOM_RESULT);
	input CLK;
	input RESET;
	input [15:0]SEED;
	output reg [15:0]RANDOM_RESULT;

	/*
	经验证，反馈系数为0111000111010110时随机循环达到最大，为65535
	*/

	always @(posedge CLK)begin
		if(RESET)begin
			RANDOM_RESULT<=SEED;
		end
		else begin
			RANDOM_RESULT[0]<=RANDOM_RESULT[15];
			RANDOM_RESULT[1]<=RANDOM_RESULT[0]^RANDOM_RESULT[15];
			RANDOM_RESULT[2]<=RANDOM_RESULT[1]^RANDOM_RESULT[15];
			RANDOM_RESULT[3]<=RANDOM_RESULT[2]^RANDOM_RESULT[15];
			RANDOM_RESULT[4]<=RANDOM_RESULT[3];
			RANDOM_RESULT[5]<=RANDOM_RESULT[4];
			RANDOM_RESULT[6]<=RANDOM_RESULT[5];
			RANDOM_RESULT[7]<=RANDOM_RESULT[6]^RANDOM_RESULT[15];
			RANDOM_RESULT[8]<=RANDOM_RESULT[7]^RANDOM_RESULT[15];
			RANDOM_RESULT[9]<=RANDOM_RESULT[8]^RANDOM_RESULT[15];
			RANDOM_RESULT[10]<=RANDOM_RESULT[9];
			RANDOM_RESULT[11]<=RANDOM_RESULT[10]^RANDOM_RESULT[15];
			RANDOM_RESULT[12]<=RANDOM_RESULT[11];
			RANDOM_RESULT[13]<=RANDOM_RESULT[12]^RANDOM_RESULT[15];
			RANDOM_RESULT[14]<=RANDOM_RESULT[13]^RANDOM_RESULT[15];
			RANDOM_RESULT[15]<=RANDOM_RESULT[14];
		end
	end
endmodule